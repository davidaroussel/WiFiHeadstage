component CLK_48MHz is
    port(
        ref_clk_i: in std_logic;
        rst_n_i: in std_logic;
        outcore_o: out std_logic;
        outglobal_o: out std_logic
    );
end component;

__: CLK_48MHz port map(
    ref_clk_i=>,
    rst_n_i=>,
    outcore_o=>,
    outglobal_o=>
);
